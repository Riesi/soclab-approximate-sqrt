--------------------------------------------------------
-- Copyright (C) 2021 Christoph Buchner under AGPLv3
--------------------------------------------------------

package Common is 
    type parity is (none,even,odd);
    type flow_ctr is (none,xon,rts,dsr);
end Common;
